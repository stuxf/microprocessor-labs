
/////////////////////////////////////////////
// sbox
//   Infamous AES byte substitutions with magic numbers
//   Synchronous version which is mapped to embedded block RAMs (EBR)
//   Section 5.1.1, Figure 7
/////////////////////////////////////////////
module sbox_sync (
    input  logic [7:0] a,
    input   logic    clk,
    output  logic [7:0] y
);

  // sbox implemented as a ROM
  // This module is synchronous and will be inferred using BRAMs (Block RAMs)
  logic [7:0] sbox[256];

  initial $readmemh("sbox.txt", sbox);

  // Synchronous version
  always_ff @(posedge clk) begin
    y <= sbox[a];
  end
endmodule
