/* 
 * Stephen Xu
 * November 4th, 2024
 * stxu@g.hmc.edu
 * This module performs SubBytes for aes
 * Applies sbox to each byte
 */
module SubBytes(
    input logic clk,
    input logic en,
    input logic[127:0] in,
    output logic[127:0] out
);

endmodule