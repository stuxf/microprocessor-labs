/* 
 * Stephen Xu
 * September 5th, 2024
 * stxu@g.hmc.edu
 * This creates a fractional clock divider
 * Uses the built in High Speed Oscillator
 */

module fractional_divider(
    input logic reset,
);

endmodule