/*
 * Stephen Xu
 * November 4th, 2024
 * stxu@g.hmc.edu
 * This module performs key expansion for aes
 * Generates round keys from key
 */
module KeyExpansion (
    input logic clk,
    input logic [127:0] inkey,
    output logic [127:0] outkey
);

  // Some sort of SubWord

endmodule
